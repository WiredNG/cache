package WiredL1Storage;

module mkWiredL1Storage();
    // 64-Bits wordsize
    // Banked data storage

    // Tag storage shared between Pipeline and manager.
endmodule

endpackage